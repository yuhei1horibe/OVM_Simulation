//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/05/2019 04:51:20 PM
// Design Name: 
// Module Name: PWM_UNIT_TEST
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`ifndef TRANS_GUARD
`define TRANS_GUARD

`include "ovm_macros.svh"
import ovm_pkg::*;

// Transaction generates patterns with constraints
// transaction is generated by generator.
class pwm_transaction extends ovm_sequence_item;
    // Define transaction pattern
    rand bit [7:0] pwm_value;
    rand bit [7:0] pwm_range;
    bit            pwm_en;

    constraint val_leq_range { pwm_value <= pwm_range; };
    constraint pwm_enable    { pwm_en    == 1'b1; };

    `ovm_object_utils_begin(pwm_transaction)
        `ovm_field_int(pwm_value, OVM_ALL_ON + OVM_DEC)
        `ovm_field_int(pwm_range, OVM_ALL_ON + OVM_DEC)
    `ovm_object_utils_end
endclass

`endif
